module test(a)

endmodule
